* C:\Users\OS1\DZ1.sch

* Schematics Version 9.1 - Web Update 1
* Fri May 14 19:18:13 2021



** Analysis setup **
.tran 1ns 500us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "dig_io.lib"
.lib "74hc.lib"
.lib "nom.lib"

.INC "DZ1.net"
.INC "DZ1.als"


.probe


.END
